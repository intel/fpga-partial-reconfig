// Copyright (c) Intel Corporation
//  
// Permission is hereby granted, free of charge, to any person obtaining a
// copy of this software and associated documentation files (the
// "Software"), to deal in the Software without restriction, including
// without limitation the rights to use, copy, modify, merge, publish,
// distribute, sublicense, and/or sell copies of the Software, and to
// permit persons to whom the Software is furnished to do so, subject to
// the following conditions:
//  
// The above copyright notice and this permission notice shall be included
// in all copies or substantial portions of the Software.
//  
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
// OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
// IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY
// CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
// TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
// SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.

module bus_pipe(clock,
		in,
		out);

   parameter WIDTH = 1;
   parameter DEPTH = 1;

   input     logic  clock;
   input     logic [WIDTH-1:0]  in;
   output    logic [WIDTH-1:0] out;

   logic [WIDTH-1:0] pipe [DEPTH-1:0] /* synthesis ramstyle = "logic" */;

   genvar 	     i;
   generate
      for (i = 0; i < DEPTH; i = i + 1) begin : block
         if (i == 0)
           always_ff @(posedge clock)
             pipe[i] <= in;
         else
           always_ff @(posedge clock)
             pipe[i] <= pipe[i-1];
      end
   endgenerate

   generate
      if (DEPTH == 0)
        assign out = in;
      else
        assign out = pipe[DEPTH-1];
   endgenerate

endmodule // bus_pipe

