`timescale 1 ps / 1 ps
`default_nettype none

// This is a template for extending the reference design to include a new persona.
// To use, define PR_CUSTOM_PERSONA in the synthesis revision qsf of your persona.

module pr_logic_template 
(
    input wire         pr_region_clk , 
    input wire         pr_logic_rst , 
    // DDR4 interface
    input wire         emif_avmm_waitrequest , 
    input wire [511:0] emif_avmm_readdata , 
    input wire         emif_avmm_readdatavalid , 
    output reg [ 4:0]  emif_avmm_burstcount , 
    output reg [511:0] emif_avmm_writedata , 
    output reg [ 30:0] emif_avmm_address , 
    output reg         emif_avmm_write , 
    output reg         emif_avmm_read , 
    output reg [ 63:0] emif_avmm_byteenable , 
    // AVMM interface
    output reg         pr_region_avmm_waitrequest , 
    output reg [ 31:0] pr_region_avmm_readdata , 
    output reg         pr_region_avmm_readdatavalid, 
    input wire [ 0:0]  pr_region_avmm_burstcount , 
    input wire [ 31:0] pr_region_avmm_writedata , 
    input wire [ 13:0] pr_region_avmm_address , 
    input wire         pr_region_avmm_write , 
    input wire         pr_region_avmm_read , 
    input wire [ 3:0]  pr_region_avmm_byteenable
    );

   //Define Number of IO registers, base case is 8 input and 8 output
   //Additional regisetrs requires modification of the reg_file.qsys
   localparam REG_FILE_IO_SIZE = 8;
   wire                clr_io_reg;

   wire [31:0]         host_pr[0:REG_FILE_IO_SIZE-1];
   wire [31:0]         pr_host [0:REG_FILE_IO_SIZE-1];

   wire [31:0]         persona_id;
   wire [31:0]         host_cntrl_register;

   `PR_CUSTOM_PERSONA #( .REG_FILE_IO_SIZE(REG_FILE_IO_SIZE) ) 
   u_pr_logic 
   (
      //clock
      .clk                       (pr_region_clk),                      
      
      //active low reset, defined by hardware
      .pr_logic_rst                     (pr_logic_rst),   
      .clr_io_reg                  (clr_io_reg),                      

      //Persona identification register, used by host in host program
      .persona_id                (persona_id),                     

      //Host control register, used for control signals.
      .host_cntrl_register       (host_cntrl_register),   

      // 8 registers for host -> PR logic communication
      .host_pr                   (host_pr),                      
      // 8 Registers for PR logic -> host communication
      .pr_host                   (pr_host),

      //DDR4 Reset
      .emif_avmm_waitrequest     (emif_avmm_waitrequest),                
      .emif_avmm_readdata        (emif_avmm_readdata),                   
      .emif_avmm_readdatavalid   (emif_avmm_readdatavalid),              
      .emif_avmm_burstcount      (emif_avmm_burstcount),                 
      .emif_avmm_writedata       (emif_avmm_writedata),                  
      .emif_avmm_address         (emif_avmm_address),                    
      .emif_avmm_write           (emif_avmm_write),                      
      .emif_avmm_read            (emif_avmm_read),                       
      .emif_avmm_byteenable      (emif_avmm_byteenable)                 
   );

   //////Register Address Map//////////////////
   //    reg_file_persona_id         = 0x0000
   //    reg_file_control_register   = 0x0010
   //    reg_file_pr_host_0          = 0x0020
   //    reg_file_pr_host_1          = 0x0030
   //    reg_file_pr_host_2          = 0x0040
   //    reg_file_pr_host_3          = 0x0050
   //    reg_file_pr_host_4          = 0x0060
   //    reg_file_pr_host_5          = 0x0070
   //    reg_file_pr_host_6          = 0x0080
   //    reg_file_pr_host_7          = 0x0090
   //    reg_file_host_pr_0          = 0x00a0
   //    reg_file_host_pr_1          = 0x00b0
   //    reg_file_host_pr_2          = 0x00c0
   //    reg_file_host_pr_3          = 0x00d0
   //    reg_file_host_pr_4          = 0x00e0
   //    reg_file_host_pr_5          = 0x00f0
   //    reg_file_host_pr_6          = 0x0100
   //    reg_file_host_pr_7          = 0x0110
   ////////////////////////////////////////////   
   reg_file u_reg_file 
      (
         //Clocking and Hardware Reset
         .reg_file_clock_clk_clk                   (pr_region_clk),
         .reg_file_hw_rst_reset                (pr_logic_rst),
         .reg_file_io_clr_reset                (clr_io_reg),
          
         //PR Identification register
         .reg_file_persona_id_export               (persona_id),

         //Host Controlled Reset
         .reg_file_control_register_export         (host_cntrl_register),

         //Avalon MM Interface
         .reg_file_mm_bridge_s0_waitrequest      (pr_region_avmm_waitrequest),
         .reg_file_mm_bridge_s0_readdata         (pr_region_avmm_readdata),
         .reg_file_mm_bridge_s0_readdatavalid    (pr_region_avmm_readdatavalid),
         .reg_file_mm_bridge_s0_burstcount       (pr_region_avmm_burstcount),
         .reg_file_mm_bridge_s0_writedata        (pr_region_avmm_writedata),
         .reg_file_mm_bridge_s0_address          (pr_region_avmm_address),
         .reg_file_mm_bridge_s0_write            (pr_region_avmm_write),
         .reg_file_mm_bridge_s0_read             (pr_region_avmm_read),
         .reg_file_mm_bridge_s0_byteenable       (pr_region_avmm_byteenable),

         //Host -> PR System registers
         .reg_file_host_pr_0_export                (host_pr[0]),
         .reg_file_host_pr_1_export                (host_pr[1]),
         .reg_file_host_pr_2_export                (host_pr[2]),
         .reg_file_host_pr_3_export                (host_pr[3]),
         .reg_file_host_pr_4_export                (host_pr[4]),
         .reg_file_host_pr_5_export                (host_pr[5]),
         .reg_file_host_pr_6_export                (host_pr[6]),
         .reg_file_host_pr_7_export                (host_pr[7]),

         // PR System -> Host registers
         .reg_file_pr_host_0_export                (pr_host[0]),
         .reg_file_pr_host_1_export                (pr_host[1]),
         .reg_file_pr_host_2_export                (pr_host[2]),
         .reg_file_pr_host_3_export                (pr_host[3]),
         .reg_file_pr_host_4_export                (pr_host[4]),
         .reg_file_pr_host_5_export                (pr_host[5]),
         .reg_file_pr_host_6_export                (pr_host[6]),
         .reg_file_pr_host_7_export                (pr_host[7])                    

      );
endmodule
