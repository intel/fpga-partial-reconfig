`ifndef INC_DESIGN_TOP_SIM_PKG_SV
`define INC_DESIGN_TOP_SIM_PKG_SV

`include "uvm_macros.svh"

package design_top_sim_pkg;
   import uvm_pkg::*;

   `include "region0_prblock_listener.sv"

   `include "sim_reporting.sv"
   `include "sb_predictor_base.sv"
   `include "sb_predictor_base.sv"
   `include "sb_predict.sv"
   `include "scoreboard.sv"
   `include "environment.sv"
   //`include "base_test.sv"

   //`include "persona_base_sequence_lib.sv"
   //`include "basic_arith_sequence_lib.sv"
   //`include "region0_pr_sequence_lib.sv"
   
endpackage


`endif //INC_DESIGN_TOP_SIM_PKG_SV
