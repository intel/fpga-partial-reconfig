// Copyright (c) Intel Corporation
//  
// Permission is hereby granted, free of charge, to any person obtaining a
// copy of this software and associated documentation files (the
// "Software"), to deal in the Software without restriction, including
// without limitation the rights to use, copy, modify, merge, publish,
// distribute, sublicense, and/or sell copies of the Software, and to
// permit persons to whom the Software is furnished to do so, subject to
// the following conditions:
//  
// The above copyright notice and this permission notice shall be included
// in all copies or substantial portions of the Software.
//  
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
// OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
// IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY
// CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
// TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
// SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.

module fifo_control(clk,
                    incr_waddr,
                    waddr,                  
                    incr_raddr,
                    raddr);

   parameter ADDR_WIDTH=5;
   
   input logic clk;
   input logic incr_waddr;
   output logic [ADDR_WIDTH-1:0] waddr;
   input logic incr_raddr;
   output logic [ADDR_WIDTH-1:0] raddr;

   always_ff @(posedge clk)
     if (incr_waddr)
       waddr <= waddr + 'b1;

   always_ff @(posedge clk)
     if (incr_raddr)
       raddr <= raddr + 'b1;
      
endmodule // fifo_control
