module sim_top();
   testbench tb();
endmodule
