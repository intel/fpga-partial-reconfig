// Copyright (c) 2001-2018 Intel Corporation
//  
// Permission is hereby granted, free of charge, to any person obtaining a
// copy of this software and associated documentation files (the
// "Software"), to deal in the Software without restriction, including
// without limitation the rights to use, copy, modify, merge, publish,
// distribute, sublicense, and/or sell copies of the Software, and to
// permit persons to whom the Software is furnished to do so, subject to
// the following conditions:
//  
// The above copyright notice and this permission notice shall be included
// in all copies or substantial portions of the Software.
//  
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
// OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
// IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY
// CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
// TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
// SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.

`ifndef INC_RESET_WATCHDOG_SV
`define INC_RESET_WATCHDOG_SV

class reset_watchdog_c extends uvm_object;

   `uvm_object_utils(reset_watchdog_c)

   virtual reset_watchdog_if vif;

   function new(string name = "reset_watchdog");
      super.new(name);
   endfunction

   task run();

      // Wait for reset complete
      `uvm_info("TST", "Waiting for reset complete", UVM_LOW)
      fork : wait_reset_complete
         begin
            while (vif.reset != 1'b0) begin
               @vif.cb1;
            end
         end
         begin
            #100000 `uvm_fatal("TST", "Reset 1 not complete")
            $finish;
         end
      join_any
      disable wait_reset_complete;
      `uvm_info("TST", "Reset 1 complete", UVM_LOW)
   
      // Post reset cycles
      repeat(10) @vif.cb1;
   
   endtask: run

endclass

`endif
